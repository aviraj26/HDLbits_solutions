module top_module(
    input clk,
    input load,
    input ena,
    input [1:0] amount,
    input [63:0] data,
    output reg [63:0] q); 
parameter lt1 = 2'b00
		 ,lt8 = 2'b01
         ,rt1 = 2'b10
		 ,rt8 = 2'b11;
    always @(posedge clk) begin
        if(load) q <= data;
        else if(ena) begin
            case(amount)
                lt1: q <= {q[62:0], 1'b0};
                lt8: q <= {q[55:0], 8'b0};
                rt1: q <= {q[63], q[63:1]};
                rt8: q <= {{8{q[63]}}, q[63:8]};
            endcase
        end    
    end
endmodule
