module top_module ( input x, input y, output z );
    xnor g(z,x,y);
endmodule
